// Copyright 2025 Google LLC
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

//----------------------------------------------------------------------------
// Description:covergroup for RV32 Zbb instruction
//----------------------------------------------------------------------------
covergroup cvgrp_RV32_Zbb;

   option.per_instance = 1;

   //base cover
   andn: coverpoint rv32zbb_trans.inst_name iff(rv32zbb_trans.trap==0) {
      bins b0 = {ANDN};
      option.weight = 1;
    }

   orn: coverpoint rv32zbb_trans.inst_name iff(rv32zbb_trans.trap==0) {
      bins b0 = {ORN};
      option.weight = 1;
    }

   xnor_: coverpoint rv32zbb_trans.inst_name iff(rv32zbb_trans.trap==0) {
      bins b0 = {XNOR};
      option.weight = 1;
    }

   clz: coverpoint rv32zbb_trans.inst_name iff(rv32zbb_trans.trap==0) {
      bins b0 = {CLZ};
      option.weight = 1;
    }

   ctz: coverpoint rv32zbb_trans.inst_name iff(rv32zbb_trans.trap==0) {
      bins b0 = {CTZ};
      option.weight = 1;
    }

   cpop: coverpoint rv32zbb_trans.inst_name iff(rv32zbb_trans.trap==0) {
      bins b0 = {CPOP};
      option.weight = 1;
    }

   max: coverpoint rv32zbb_trans.inst_name iff(rv32zbb_trans.trap==0) {
      bins b0 = {MAX};
      option.weight = 1;
    }

   maxu: coverpoint rv32zbb_trans.inst_name iff(rv32zbb_trans.trap==0) {
      bins b0 = {MAXU};
      option.weight = 1;
    }

   min: coverpoint rv32zbb_trans.inst_name iff(rv32zbb_trans.trap==0) {
      bins b0 = {MIN};
      option.weight = 1;
    }

   minu: coverpoint rv32zbb_trans.inst_name iff(rv32zbb_trans.trap==0) {
      bins b0 = {MINU};
      option.weight = 1;
    }

   sext_b: coverpoint rv32zbb_trans.inst_name iff(rv32zbb_trans.trap==0) {
      bins b0 = {SEXT_B};
      option.weight = 1;
    }

   sext_h: coverpoint rv32zbb_trans.inst_name iff(rv32zbb_trans.trap==0) {
      bins b0 = {SEXT_H};
      option.weight = 1;
    }

   zext_h: coverpoint rv32zbb_trans.inst_name iff(rv32zbb_trans.trap==0) {
      bins b0 = {ZEXT_H};
      option.weight = 1;
    }

   rol: coverpoint rv32zbb_trans.inst_name iff(rv32zbb_trans.trap==0) {
      bins b0 = {ROL};
      option.weight = 1;
    }

   ror: coverpoint rv32zbb_trans.inst_name iff(rv32zbb_trans.trap==0) {
      bins b0 = {ROR};
      option.weight = 1;
    }

   rori: coverpoint rv32zbb_trans.inst_name iff(rv32zbb_trans.trap==0) {
      bins b0 = {RORI};
      option.weight = 1;
    }

   orc_b: coverpoint rv32zbb_trans.inst_name iff(rv32zbb_trans.trap==0) {
      bins b0 = {ORC_B};
      option.weight = 1;
    }

   rev8: coverpoint rv32zbb_trans.inst_name iff(rv32zbb_trans.trap==0) {
      bins b0 = {REV8};
      option.weight = 1;
    }

   //RD (GPR) register assignment,x0 always 0
   rd_addr: coverpoint rv32zbb_trans.rd_addr iff(rv32zbb_trans.trap==0) {
      bins b0 = {0};
      bins b1 = {1};
      bins b2 = {2};
      bins b3 = {3};
      bins b4 = {4};
      bins b5 = {5};
      bins b6 = {6};
      bins b7 = {7};
      bins b8 = {8};
      bins b9 = {9};
      bins b10 = {10};
      bins b11 = {11};
      bins b12 = {12};
      bins b13 = {13};
      bins b14 = {14};
      bins b15 = {15};
      bins b16 = {16};
      bins b17 = {17};
      bins b18 = {18};
      bins b19 = {19};
      bins b20 = {20};
      bins b21 = {21};
      bins b22 = {22};
      bins b23 = {23};
      bins b24 = {24};
      bins b25 = {25};
      bins b26 = {26};
      bins b27 = {27};
      bins b28 = {28};
      bins b29 = {29};
      bins b30 = {30};
      bins b31 = {31};
      option.weight = 1;
    }

   //RS1 (GPR) register assignment
   rs1_addr: coverpoint rv32zbb_trans.rs1_addr iff(rv32zbb_trans.trap==0) {
      bins b0 = {0};
      bins b1 = {1};
      bins b2 = {2};
      bins b3 = {3};
      bins b4 = {4};
      bins b5 = {5};
      bins b6 = {6};
      bins b7 = {7};
      bins b8 = {8};
      bins b9 = {9};
      bins b10 = {10};
      bins b11 = {11};
      bins b12 = {12};
      bins b13 = {13};
      bins b14 = {14};
      bins b15 = {15};
      bins b16 = {16};
      bins b17 = {17};
      bins b18 = {18};
      bins b19 = {19};
      bins b20 = {20};
      bins b21 = {21};
      bins b22 = {22};
      bins b23 = {23};
      bins b24 = {24};
      bins b25 = {25};
      bins b26 = {26};
      bins b27 = {27};
      bins b28 = {28};
      bins b29 = {29};
      bins b30 = {30};
      bins b31 = {31};
      option.weight = 1;
    }

   //RS2 (GPR) register assignment
   rs2_addr: coverpoint rv32zbb_trans.rs2_addr iff(rv32zbb_trans.trap==0) {
      bins b0 = {0};
      bins b1 = {1};
      bins b2 = {2};
      bins b3 = {3};
      bins b4 = {4};
      bins b5 = {5};
      bins b6 = {6};
      bins b7 = {7};
      bins b8 = {8};
      bins b9 = {9};
      bins b10 = {10};
      bins b11 = {11};
      bins b12 = {12};
      bins b13 = {13};
      bins b14 = {14};
      bins b15 = {15};
      bins b16 = {16};
      bins b17 = {17};
      bins b18 = {18};
      bins b19 = {19};
      bins b20 = {20};
      bins b21 = {21};
      bins b22 = {22};
      bins b23 = {23};
      bins b24 = {24};
      bins b25 = {25};
      bins b26 = {26};
      bins b27 = {27};
      bins b28 = {28};
      bins b29 = {29};
      bins b30 = {30};
      bins b31 = {31};
      option.weight = 1;
    }

   //shamt toggle bits
   shamt_val: coverpoint unsigned'(rv32zbb_trans.shamt) iff(rv32zbb_trans.inst_name==coralnpu_rvvi_agent_pkg::RORI&&rv32zbb_trans.trap==0) {
      wildcard bins b_1_0_0    = (5'b????1=>5'b????0);
      wildcard bins b_1_0_1    = (5'b???1?=>5'b???0?);
      wildcard bins b_1_0_2    = (5'b??1??=>5'b??0??);
      wildcard bins b_1_0_3    = (5'b?1???=>5'b?0???);
      wildcard bins b_1_0_4    = (5'b1????=>5'b0????);
      wildcard bins b_0_1_0    = (5'b????0=>5'b????1);
      wildcard bins b_0_1_1    = (5'b???0?=>5'b???1?);
      wildcard bins b_0_1_2    = (5'b??0??=>5'b??1??);
      wildcard bins b_0_1_3    = (5'b?0???=>5'b?1???);
      wildcard bins b_0_1_4    = (5'b0????=>5'b1????);
      option.weight = 1;
    }

   //shamt special values
   shamt_sp_val: coverpoint unsigned'(rv32zbb_trans.shamt) iff(rv32zbb_trans.inst_name==coralnpu_rvvi_agent_pkg::RORI&&rv32zbb_trans.trap==0) {
      bins b0 = {5'b0};
      bins b1 = {5'b00001};
      bins b2 = {5'b11111};
      bins b3 = {5'b10000};
      bins b4 = {5'b10001};
      option.weight = 1;
    }

   //shamt special values
   rd_val: coverpoint unsigned'(rv32zbb_trans.rd_val) iff(rv32zbb_trans.trap==0) {
      wildcard bins b_1_0_0    = (32'b???????????????????????????????1=>32'b???????????????????????????????0);
      wildcard bins b_1_0_1    = (32'b??????????????????????????????1?=>32'b??????????????????????????????0?);
      wildcard bins b_1_0_2    = (32'b?????????????????????????????1??=>32'b?????????????????????????????0??);
      wildcard bins b_1_0_3    = (32'b????????????????????????????1???=>32'b????????????????????????????0???);
      wildcard bins b_1_0_4    = (32'b???????????????????????????1????=>32'b???????????????????????????0????);
      wildcard bins b_1_0_5    = (32'b??????????????????????????1?????=>32'b??????????????????????????0?????);
      wildcard bins b_1_0_6    = (32'b?????????????????????????1??????=>32'b?????????????????????????0??????);
      wildcard bins b_1_0_7    = (32'b????????????????????????1???????=>32'b????????????????????????0???????);
      wildcard bins b_1_0_8    = (32'b???????????????????????1????????=>32'b???????????????????????0????????);
      wildcard bins b_1_0_9    = (32'b??????????????????????1?????????=>32'b??????????????????????0?????????);
      wildcard bins b_1_0_10    = (32'b?????????????????????1??????????=>32'b?????????????????????0??????????);
      wildcard bins b_1_0_11    = (32'b????????????????????1???????????=>32'b????????????????????0???????????);
      wildcard bins b_1_0_12    = (32'b???????????????????1????????????=>32'b???????????????????0????????????);
      wildcard bins b_1_0_13    = (32'b??????????????????1?????????????=>32'b??????????????????0?????????????);
      wildcard bins b_1_0_14    = (32'b?????????????????1??????????????=>32'b?????????????????0??????????????);
      wildcard bins b_1_0_15    = (32'b????????????????1???????????????=>32'b????????????????0???????????????);
      wildcard bins b_1_0_16    = (32'b???????????????1????????????????=>32'b???????????????0????????????????);
      wildcard bins b_1_0_17    = (32'b??????????????1?????????????????=>32'b??????????????0?????????????????);
      wildcard bins b_1_0_18    = (32'b?????????????1??????????????????=>32'b?????????????0??????????????????);
      wildcard bins b_1_0_19    = (32'b????????????1???????????????????=>32'b????????????0???????????????????);
      wildcard bins b_1_0_20    = (32'b???????????1????????????????????=>32'b???????????0????????????????????);
      wildcard bins b_1_0_21    = (32'b??????????1?????????????????????=>32'b??????????0?????????????????????);
      wildcard bins b_1_0_22    = (32'b?????????1??????????????????????=>32'b?????????0??????????????????????);
      wildcard bins b_1_0_23    = (32'b????????1???????????????????????=>32'b????????0???????????????????????);
      wildcard bins b_1_0_24    = (32'b???????1????????????????????????=>32'b???????0????????????????????????);
      wildcard bins b_1_0_25    = (32'b??????1?????????????????????????=>32'b??????0?????????????????????????);
      wildcard bins b_1_0_26    = (32'b?????1??????????????????????????=>32'b?????0??????????????????????????);
      wildcard bins b_1_0_27    = (32'b????1???????????????????????????=>32'b????0???????????????????????????);
      wildcard bins b_1_0_28    = (32'b???1????????????????????????????=>32'b???0????????????????????????????);
      wildcard bins b_1_0_29    = (32'b??1?????????????????????????????=>32'b??0?????????????????????????????);
      wildcard bins b_1_0_30    = (32'b?1??????????????????????????????=>32'b?0??????????????????????????????);
      wildcard bins b_1_0_31    = (32'b1???????????????????????????????=>32'b0???????????????????????????????);
      wildcard bins b_0_1_0    = (32'b???????????????????????????????0=>32'b???????????????????????????????1);
      wildcard bins b_0_1_1    = (32'b??????????????????????????????0?=>32'b??????????????????????????????1?);
      wildcard bins b_0_1_2    = (32'b?????????????????????????????0??=>32'b?????????????????????????????1??);
      wildcard bins b_0_1_3    = (32'b????????????????????????????0???=>32'b????????????????????????????1???);
      wildcard bins b_0_1_4    = (32'b???????????????????????????0????=>32'b???????????????????????????1????);
      wildcard bins b_0_1_5    = (32'b??????????????????????????0?????=>32'b??????????????????????????1?????);
      wildcard bins b_0_1_6    = (32'b?????????????????????????0??????=>32'b?????????????????????????1??????);
      wildcard bins b_0_1_7    = (32'b????????????????????????0???????=>32'b????????????????????????1???????);
      wildcard bins b_0_1_8    = (32'b???????????????????????0????????=>32'b???????????????????????1????????);
      wildcard bins b_0_1_9    = (32'b??????????????????????0?????????=>32'b??????????????????????1?????????);
      wildcard bins b_0_1_10    = (32'b?????????????????????0??????????=>32'b?????????????????????1??????????);
      wildcard bins b_0_1_11    = (32'b????????????????????0???????????=>32'b????????????????????1???????????);
      wildcard bins b_0_1_12    = (32'b???????????????????0????????????=>32'b???????????????????1????????????);
      wildcard bins b_0_1_13    = (32'b??????????????????0?????????????=>32'b??????????????????1?????????????);
      wildcard bins b_0_1_14    = (32'b?????????????????0??????????????=>32'b?????????????????1??????????????);
      wildcard bins b_0_1_15    = (32'b????????????????0???????????????=>32'b????????????????1???????????????);
      wildcard bins b_0_1_16    = (32'b???????????????0????????????????=>32'b???????????????1????????????????);
      wildcard bins b_0_1_17    = (32'b??????????????0?????????????????=>32'b??????????????1?????????????????);
      wildcard bins b_0_1_18    = (32'b?????????????0??????????????????=>32'b?????????????1??????????????????);
      wildcard bins b_0_1_19    = (32'b????????????0???????????????????=>32'b????????????1???????????????????);
      wildcard bins b_0_1_20    = (32'b???????????0????????????????????=>32'b???????????1????????????????????);
      wildcard bins b_0_1_21    = (32'b??????????0?????????????????????=>32'b??????????1?????????????????????);
      wildcard bins b_0_1_22    = (32'b?????????0??????????????????????=>32'b?????????1??????????????????????);
      wildcard bins b_0_1_23    = (32'b????????0???????????????????????=>32'b????????1???????????????????????);
      wildcard bins b_0_1_24    = (32'b???????0????????????????????????=>32'b???????1????????????????????????);
      wildcard bins b_0_1_25    = (32'b??????0?????????????????????????=>32'b??????1?????????????????????????);
      wildcard bins b_0_1_26    = (32'b?????0??????????????????????????=>32'b?????1??????????????????????????);
      wildcard bins b_0_1_27    = (32'b????0???????????????????????????=>32'b????1???????????????????????????);
      wildcard bins b_0_1_28    = (32'b???0????????????????????????????=>32'b???1????????????????????????????);
      wildcard bins b_0_1_29    = (32'b??0?????????????????????????????=>32'b??1?????????????????????????????);
      wildcard bins b_0_1_30    = (32'b?0??????????????????????????????=>32'b?1??????????????????????????????);
      wildcard bins b_0_1_31    = (32'b0???????????????????????????????=>32'b1???????????????????????????????);
      option.weight = 1;
    }

   //RD special values
   rd_sp_val: coverpoint unsigned'(rv32zbb_trans.rd_val) iff(rv32zbb_trans.trap==0) {
      bins b0 = {32'b0};
      bins b1 = {32'b00000000000000000000000000000001};
      bins b2 = {32'b11111111111111111111111111111111};
      bins b3 = {32'b01111111111111111111111111111111};
      bins b4 = {32'b10000000000000000000000000000000};
      bins b5 = {32'b10000000000000000000000000000001};
      option.weight = 1;
    }

   //RD value sign
   rd_val_sign: coverpoint rv32zbb_trans.rd_val iff(rv32zbb_trans.trap==0) {
      bins b0 = {[$:-1]};
      bins b1 = {[1:$]};
      option.weight = 1;
    }

   //RS1 toggle bits
   rs1_val: coverpoint unsigned'(rv32zbb_trans.rs1_val) iff(rv32zbb_trans.trap==0) {
      wildcard bins b_1_0_0    = (32'b???????????????????????????????1=>32'b???????????????????????????????0);
      wildcard bins b_1_0_1    = (32'b??????????????????????????????1?=>32'b??????????????????????????????0?);
      wildcard bins b_1_0_2    = (32'b?????????????????????????????1??=>32'b?????????????????????????????0??);
      wildcard bins b_1_0_3    = (32'b????????????????????????????1???=>32'b????????????????????????????0???);
      wildcard bins b_1_0_4    = (32'b???????????????????????????1????=>32'b???????????????????????????0????);
      wildcard bins b_1_0_5    = (32'b??????????????????????????1?????=>32'b??????????????????????????0?????);
      wildcard bins b_1_0_6    = (32'b?????????????????????????1??????=>32'b?????????????????????????0??????);
      wildcard bins b_1_0_7    = (32'b????????????????????????1???????=>32'b????????????????????????0???????);
      wildcard bins b_1_0_8    = (32'b???????????????????????1????????=>32'b???????????????????????0????????);
      wildcard bins b_1_0_9    = (32'b??????????????????????1?????????=>32'b??????????????????????0?????????);
      wildcard bins b_1_0_10    = (32'b?????????????????????1??????????=>32'b?????????????????????0??????????);
      wildcard bins b_1_0_11    = (32'b????????????????????1???????????=>32'b????????????????????0???????????);
      wildcard bins b_1_0_12    = (32'b???????????????????1????????????=>32'b???????????????????0????????????);
      wildcard bins b_1_0_13    = (32'b??????????????????1?????????????=>32'b??????????????????0?????????????);
      wildcard bins b_1_0_14    = (32'b?????????????????1??????????????=>32'b?????????????????0??????????????);
      wildcard bins b_1_0_15    = (32'b????????????????1???????????????=>32'b????????????????0???????????????);
      wildcard bins b_1_0_16    = (32'b???????????????1????????????????=>32'b???????????????0????????????????);
      wildcard bins b_1_0_17    = (32'b??????????????1?????????????????=>32'b??????????????0?????????????????);
      wildcard bins b_1_0_18    = (32'b?????????????1??????????????????=>32'b?????????????0??????????????????);
      wildcard bins b_1_0_19    = (32'b????????????1???????????????????=>32'b????????????0???????????????????);
      wildcard bins b_1_0_20    = (32'b???????????1????????????????????=>32'b???????????0????????????????????);
      wildcard bins b_1_0_21    = (32'b??????????1?????????????????????=>32'b??????????0?????????????????????);
      wildcard bins b_1_0_22    = (32'b?????????1??????????????????????=>32'b?????????0??????????????????????);
      wildcard bins b_1_0_23    = (32'b????????1???????????????????????=>32'b????????0???????????????????????);
      wildcard bins b_1_0_24    = (32'b???????1????????????????????????=>32'b???????0????????????????????????);
      wildcard bins b_1_0_25    = (32'b??????1?????????????????????????=>32'b??????0?????????????????????????);
      wildcard bins b_1_0_26    = (32'b?????1??????????????????????????=>32'b?????0??????????????????????????);
      wildcard bins b_1_0_27    = (32'b????1???????????????????????????=>32'b????0???????????????????????????);
      wildcard bins b_1_0_28    = (32'b???1????????????????????????????=>32'b???0????????????????????????????);
      wildcard bins b_1_0_29    = (32'b??1?????????????????????????????=>32'b??0?????????????????????????????);
      wildcard bins b_1_0_30    = (32'b?1??????????????????????????????=>32'b?0??????????????????????????????);
      wildcard bins b_1_0_31    = (32'b1???????????????????????????????=>32'b0???????????????????????????????);
      wildcard bins b_0_1_0    = (32'b???????????????????????????????0=>32'b???????????????????????????????1);
      wildcard bins b_0_1_1    = (32'b??????????????????????????????0?=>32'b??????????????????????????????1?);
      wildcard bins b_0_1_2    = (32'b?????????????????????????????0??=>32'b?????????????????????????????1??);
      wildcard bins b_0_1_3    = (32'b????????????????????????????0???=>32'b????????????????????????????1???);
      wildcard bins b_0_1_4    = (32'b???????????????????????????0????=>32'b???????????????????????????1????);
      wildcard bins b_0_1_5    = (32'b??????????????????????????0?????=>32'b??????????????????????????1?????);
      wildcard bins b_0_1_6    = (32'b?????????????????????????0??????=>32'b?????????????????????????1??????);
      wildcard bins b_0_1_7    = (32'b????????????????????????0???????=>32'b????????????????????????1???????);
      wildcard bins b_0_1_8    = (32'b???????????????????????0????????=>32'b???????????????????????1????????);
      wildcard bins b_0_1_9    = (32'b??????????????????????0?????????=>32'b??????????????????????1?????????);
      wildcard bins b_0_1_10    = (32'b?????????????????????0??????????=>32'b?????????????????????1??????????);
      wildcard bins b_0_1_11    = (32'b????????????????????0???????????=>32'b????????????????????1???????????);
      wildcard bins b_0_1_12    = (32'b???????????????????0????????????=>32'b???????????????????1????????????);
      wildcard bins b_0_1_13    = (32'b??????????????????0?????????????=>32'b??????????????????1?????????????);
      wildcard bins b_0_1_14    = (32'b?????????????????0??????????????=>32'b?????????????????1??????????????);
      wildcard bins b_0_1_15    = (32'b????????????????0???????????????=>32'b????????????????1???????????????);
      wildcard bins b_0_1_16    = (32'b???????????????0????????????????=>32'b???????????????1????????????????);
      wildcard bins b_0_1_17    = (32'b??????????????0?????????????????=>32'b??????????????1?????????????????);
      wildcard bins b_0_1_18    = (32'b?????????????0??????????????????=>32'b?????????????1??????????????????);
      wildcard bins b_0_1_19    = (32'b????????????0???????????????????=>32'b????????????1???????????????????);
      wildcard bins b_0_1_20    = (32'b???????????0????????????????????=>32'b???????????1????????????????????);
      wildcard bins b_0_1_21    = (32'b??????????0?????????????????????=>32'b??????????1?????????????????????);
      wildcard bins b_0_1_22    = (32'b?????????0??????????????????????=>32'b?????????1??????????????????????);
      wildcard bins b_0_1_23    = (32'b????????0???????????????????????=>32'b????????1???????????????????????);
      wildcard bins b_0_1_24    = (32'b???????0????????????????????????=>32'b???????1????????????????????????);
      wildcard bins b_0_1_25    = (32'b??????0?????????????????????????=>32'b??????1?????????????????????????);
      wildcard bins b_0_1_26    = (32'b?????0??????????????????????????=>32'b?????1??????????????????????????);
      wildcard bins b_0_1_27    = (32'b????0???????????????????????????=>32'b????1???????????????????????????);
      wildcard bins b_0_1_28    = (32'b???0????????????????????????????=>32'b???1????????????????????????????);
      wildcard bins b_0_1_29    = (32'b??0?????????????????????????????=>32'b??1?????????????????????????????);
      wildcard bins b_0_1_30    = (32'b?0??????????????????????????????=>32'b?1??????????????????????????????);
      wildcard bins b_0_1_31    = (32'b0???????????????????????????????=>32'b1???????????????????????????????);
      option.weight = 1;
    }

   //RS1 special values
   rs1_sp_val: coverpoint unsigned'(rv32zbb_trans.rs1_val) iff(rv32zbb_trans.trap==0) {
      bins b0 = {32'b0};
      bins b1 = {32'b00000000000000000000000000000001};
      bins b2 = {32'b11111111111111111111111111111111};
      bins b3 = {32'b01111111111111111111111111111111};
      bins b4 = {32'b10000000000000000000000000000000};
      bins b5 = {32'b10000000000000000000000000000001};
      option.weight = 1;
    }

   //RS1 value sign
   rs1_val_sign: coverpoint rv32zbb_trans.rs1_val iff(rv32zbb_trans.trap==0) {
      bins b0 = {[$:-1]};
      bins b1 = {[1:$]};
      option.weight = 1;
    }

   //RS2 toggle bits
   rs2_val: coverpoint unsigned'(rv32zbb_trans.rs2_val) iff(rv32zbb_trans.trap==0) {
      wildcard bins b_1_0_0    = (32'b???????????????????????????????1=>32'b???????????????????????????????0);
      wildcard bins b_1_0_1    = (32'b??????????????????????????????1?=>32'b??????????????????????????????0?);
      wildcard bins b_1_0_2    = (32'b?????????????????????????????1??=>32'b?????????????????????????????0??);
      wildcard bins b_1_0_3    = (32'b????????????????????????????1???=>32'b????????????????????????????0???);
      wildcard bins b_1_0_4    = (32'b???????????????????????????1????=>32'b???????????????????????????0????);
      wildcard bins b_1_0_5    = (32'b??????????????????????????1?????=>32'b??????????????????????????0?????);
      wildcard bins b_1_0_6    = (32'b?????????????????????????1??????=>32'b?????????????????????????0??????);
      wildcard bins b_1_0_7    = (32'b????????????????????????1???????=>32'b????????????????????????0???????);
      wildcard bins b_1_0_8    = (32'b???????????????????????1????????=>32'b???????????????????????0????????);
      wildcard bins b_1_0_9    = (32'b??????????????????????1?????????=>32'b??????????????????????0?????????);
      wildcard bins b_1_0_10    = (32'b?????????????????????1??????????=>32'b?????????????????????0??????????);
      wildcard bins b_1_0_11    = (32'b????????????????????1???????????=>32'b????????????????????0???????????);
      wildcard bins b_1_0_12    = (32'b???????????????????1????????????=>32'b???????????????????0????????????);
      wildcard bins b_1_0_13    = (32'b??????????????????1?????????????=>32'b??????????????????0?????????????);
      wildcard bins b_1_0_14    = (32'b?????????????????1??????????????=>32'b?????????????????0??????????????);
      wildcard bins b_1_0_15    = (32'b????????????????1???????????????=>32'b????????????????0???????????????);
      wildcard bins b_1_0_16    = (32'b???????????????1????????????????=>32'b???????????????0????????????????);
      wildcard bins b_1_0_17    = (32'b??????????????1?????????????????=>32'b??????????????0?????????????????);
      wildcard bins b_1_0_18    = (32'b?????????????1??????????????????=>32'b?????????????0??????????????????);
      wildcard bins b_1_0_19    = (32'b????????????1???????????????????=>32'b????????????0???????????????????);
      wildcard bins b_1_0_20    = (32'b???????????1????????????????????=>32'b???????????0????????????????????);
      wildcard bins b_1_0_21    = (32'b??????????1?????????????????????=>32'b??????????0?????????????????????);
      wildcard bins b_1_0_22    = (32'b?????????1??????????????????????=>32'b?????????0??????????????????????);
      wildcard bins b_1_0_23    = (32'b????????1???????????????????????=>32'b????????0???????????????????????);
      wildcard bins b_1_0_24    = (32'b???????1????????????????????????=>32'b???????0????????????????????????);
      wildcard bins b_1_0_25    = (32'b??????1?????????????????????????=>32'b??????0?????????????????????????);
      wildcard bins b_1_0_26    = (32'b?????1??????????????????????????=>32'b?????0??????????????????????????);
      wildcard bins b_1_0_27    = (32'b????1???????????????????????????=>32'b????0???????????????????????????);
      wildcard bins b_1_0_28    = (32'b???1????????????????????????????=>32'b???0????????????????????????????);
      wildcard bins b_1_0_29    = (32'b??1?????????????????????????????=>32'b??0?????????????????????????????);
      wildcard bins b_1_0_30    = (32'b?1??????????????????????????????=>32'b?0??????????????????????????????);
      wildcard bins b_1_0_31    = (32'b1???????????????????????????????=>32'b0???????????????????????????????);
      wildcard bins b_0_1_0    = (32'b???????????????????????????????0=>32'b???????????????????????????????1);
      wildcard bins b_0_1_1    = (32'b??????????????????????????????0?=>32'b??????????????????????????????1?);
      wildcard bins b_0_1_2    = (32'b?????????????????????????????0??=>32'b?????????????????????????????1??);
      wildcard bins b_0_1_3    = (32'b????????????????????????????0???=>32'b????????????????????????????1???);
      wildcard bins b_0_1_4    = (32'b???????????????????????????0????=>32'b???????????????????????????1????);
      wildcard bins b_0_1_5    = (32'b??????????????????????????0?????=>32'b??????????????????????????1?????);
      wildcard bins b_0_1_6    = (32'b?????????????????????????0??????=>32'b?????????????????????????1??????);
      wildcard bins b_0_1_7    = (32'b????????????????????????0???????=>32'b????????????????????????1???????);
      wildcard bins b_0_1_8    = (32'b???????????????????????0????????=>32'b???????????????????????1????????);
      wildcard bins b_0_1_9    = (32'b??????????????????????0?????????=>32'b??????????????????????1?????????);
      wildcard bins b_0_1_10    = (32'b?????????????????????0??????????=>32'b?????????????????????1??????????);
      wildcard bins b_0_1_11    = (32'b????????????????????0???????????=>32'b????????????????????1???????????);
      wildcard bins b_0_1_12    = (32'b???????????????????0????????????=>32'b???????????????????1????????????);
      wildcard bins b_0_1_13    = (32'b??????????????????0?????????????=>32'b??????????????????1?????????????);
      wildcard bins b_0_1_14    = (32'b?????????????????0??????????????=>32'b?????????????????1??????????????);
      wildcard bins b_0_1_15    = (32'b????????????????0???????????????=>32'b????????????????1???????????????);
      wildcard bins b_0_1_16    = (32'b???????????????0????????????????=>32'b???????????????1????????????????);
      wildcard bins b_0_1_17    = (32'b??????????????0?????????????????=>32'b??????????????1?????????????????);
      wildcard bins b_0_1_18    = (32'b?????????????0??????????????????=>32'b?????????????1??????????????????);
      wildcard bins b_0_1_19    = (32'b????????????0???????????????????=>32'b????????????1???????????????????);
      wildcard bins b_0_1_20    = (32'b???????????0????????????????????=>32'b???????????1????????????????????);
      wildcard bins b_0_1_21    = (32'b??????????0?????????????????????=>32'b??????????1?????????????????????);
      wildcard bins b_0_1_22    = (32'b?????????0??????????????????????=>32'b?????????1??????????????????????);
      wildcard bins b_0_1_23    = (32'b????????0???????????????????????=>32'b????????1???????????????????????);
      wildcard bins b_0_1_24    = (32'b???????0????????????????????????=>32'b???????1????????????????????????);
      wildcard bins b_0_1_25    = (32'b??????0?????????????????????????=>32'b??????1?????????????????????????);
      wildcard bins b_0_1_26    = (32'b?????0??????????????????????????=>32'b?????1??????????????????????????);
      wildcard bins b_0_1_27    = (32'b????0???????????????????????????=>32'b????1???????????????????????????);
      wildcard bins b_0_1_28    = (32'b???0????????????????????????????=>32'b???1????????????????????????????);
      wildcard bins b_0_1_29    = (32'b??0?????????????????????????????=>32'b??1?????????????????????????????);
      wildcard bins b_0_1_30    = (32'b?0??????????????????????????????=>32'b?1??????????????????????????????);
      wildcard bins b_0_1_31    = (32'b0???????????????????????????????=>32'b1???????????????????????????????);
      option.weight = 1;
    }

   //RS2 special values
   rs2_sp_val: coverpoint unsigned'(rv32zbb_trans.rs2_val) iff(rv32zbb_trans.trap==0) {
      bins b0 = {32'b0};
      bins b1 = {32'b00000000000000000000000000000001};
      bins b2 = {32'b11111111111111111111111111111111};
      bins b3 = {32'b01111111111111111111111111111111};
      bins b4 = {32'b10000000000000000000000000000000};
      bins b5 = {32'b10000000000000000000000000000001};
      option.weight = 1;
    }

   //RS2 value sign
   rs2_val_sign: coverpoint rv32zbb_trans.rs2_val iff(rv32zbb_trans.trap==0) {
      bins b0 = {[$:-1]};
      bins b1 = {[1:$]};
      option.weight = 1;
    }

   //war_hazard
   war_hazard_hit: coverpoint rv32zbb_trans.war_hazard_hit iff(rv32zbb_trans.trap==0) {
      bins b0 = {1};
      option.weight = 1;
    }

   //waw_hazard
   waw_hazard_hit: coverpoint rv32zbb_trans.waw_hazard_hit iff(rv32zbb_trans.trap==0) {
      bins b0 = {1};
      option.weight = 1;
    }

   //raw_hazard
   raw_hazard_hit: coverpoint rv32zbb_trans.raw_hazard_hit iff(rv32zbb_trans.trap==0) {
      bins b0 = {1};
      option.weight = 1;
    }

   // base cross
   //ANDN instruction crosspoints
   //Cross ANDN instruction and register assignment
   cr_andn_rs1_rs2_rd: cross andn,rs1_addr,rs2_addr,rd_addr {
      option.weight = 1;
   }

   //Cross ANDN instruction and RS1 toggle bits
   cr_andn_rs1_val: cross andn,rs1_val {
      option.weight = 1;
   }

   //Cross ANDN instruction and RS1 special values
   cr_andn_rs1_sp_val: cross andn,rs1_sp_val {
      option.weight = 1;
   }

   //Cross ANDN instruction and RS2 toggle bits
   cr_andn_rs2_val: cross andn,rs2_val {
      option.weight = 1;
   }

   //Cross ANDN instruction and RS2 special values
   cr_andn_rs2_sp_val: cross andn,rs2_sp_val {
      option.weight = 1;
   }

   //Cross ANDN instruction and RD toggle bits
   cr_andn_rd_val: cross andn,rd_val {
      option.weight = 1;
   }

   //Cross ANDN instruction and RD special values
   cr_andn_rd_sp_val: cross andn,rd_sp_val {
      option.weight = 1;
   }

   //Cross ANDN instruction and WAR hazard
   cr_andn_war_hazard: cross andn,war_hazard_hit {
      option.weight = 1;
   }

   //Cross ANDN instruction and WAW hazard
   cr_andn_waw_hazard: cross andn,waw_hazard_hit {
      option.weight = 1;
   }

   //Cross ANDN instruction and RAW hazard
   cr_andn_raw_hazard: cross andn,raw_hazard_hit {
      option.weight = 1;
   }

   //ORN instruction crosspoints
   //Cross ORN instruction and register assignment
   cr_orn_rs1_rs2_rd: cross orn,rs1_addr,rs2_addr,rd_addr {
      option.weight = 1;
   }

   //Cross ORN instruction and RS1 toggle bits
   cr_orn_rs1_val: cross orn,rs1_val {
      option.weight = 1;
   }

   //Cross ORN instruction and RS1 special values
   cr_orn_rs1_sp_val: cross orn,rs1_sp_val {
      option.weight = 1;
   }

   //Cross ORN instruction and RS2 toggle bits
   cr_orn_rs2_val: cross orn,rs2_val {
      option.weight = 1;
   }

   //Cross ORN instruction and RS2 special values
   cr_orn_rs2_sp_val: cross orn,rs2_sp_val {
      option.weight = 1;
   }

   //Cross ORN instruction and RD toggle bits
   cr_orn_rd_val: cross orn,rd_val {
      option.weight = 1;
   }

   //Cross ORN instruction and RD special values
   cr_orn_rd_sp_val: cross orn,rd_sp_val {
      option.weight = 1;
   }

   //Cross ORN instruction and WAR hazard
   cr_orn_war_hazard: cross orn,war_hazard_hit {
      option.weight = 1;
   }

   //Cross ORN instruction and WAW hazard
   cr_orn_waw_hazard: cross orn,waw_hazard_hit {
      option.weight = 1;
   }

   //Cross ORN instruction and RAW hazard
   cr_orn_raw_hazard: cross orn,raw_hazard_hit {
      option.weight = 1;
   }

   //XNOR instruction crosspoints
   //Cross XNOR instruction and register assignment
   cr_xnor_rs1_rs2_rd: cross xnor_,rs1_addr,rs2_addr,rd_addr {
      option.weight = 1;
   }

   //Cross XNOR instruction and RS1 toggle bits
   cr_xnor_rs1_val: cross xnor_,rs1_val {
      option.weight = 1;
   }

   //Cross XNOR instruction and RS1 special values
   cr_xnor_rs1_sp_val: cross xnor_,rs1_sp_val {
      option.weight = 1;
   }

   //Cross XNOR instruction and RS2 toggle bits
   cr_xnor_rs2_val: cross xnor_,rs2_val {
      option.weight = 1;
   }

   //Cross XNOR instruction and RS2 special values
   cr_xnor_rs2_sp_val: cross xnor_,rs2_sp_val {
      option.weight = 1;
   }

   //Cross XNOR instruction and RD toggle bits
   cr_xnor_rd_val: cross xnor_,rd_val {
      option.weight = 1;
   }

   //Cross XNOR instruction and RD special values
   cr_xnor_rd_sp_val: cross xnor_,rd_sp_val {
      option.weight = 1;
   }

   //Cross XNOR instruction and WAR hazard
   cr_xnor_war_hazard: cross xnor_,war_hazard_hit {
      option.weight = 1;
   }

   //Cross XNOR instruction and WAW hazard
   cr_xnor_waw_hazard: cross xnor_,waw_hazard_hit {
      option.weight = 1;
   }

   //Cross XNOR instruction and RAW hazard
   cr_xnor_raw_hazard: cross xnor_,raw_hazard_hit {
      option.weight = 1;
   }

   //CLZ instruction crosspoints
   //Cross CLZ instruction and register assignment
   cr_clz_rs1_rd: cross clz,rs1_addr,rd_addr {
      option.weight = 1;
   }

   //Cross CLZ instruction and RS1 toggle bits
   cr_clz_rs1_val: cross clz,rs1_val {
      option.weight = 1;
   }

   //Cross CLZ instruction and RS1 special values
   cr_clz_rs1_sp_val: cross clz,rs1_sp_val {
      option.weight = 1;
   }

   //Cross CLZ instruction and RD toggle bits
   cr_clz_rd_val: cross clz,rd_val {
      option.weight = 1;
   }

   //Cross CLZ instruction and RD special values
   cr_clz_rd_sp_val: cross clz,rd_sp_val {
      option.weight = 1;
   }

   //Cross CLZ instruction and WAR hazard
   cr_clz_war_hazard: cross clz,war_hazard_hit {
      option.weight = 1;
   }

   //Cross CLZ instruction and WAW hazard
   cr_clz_waw_hazard: cross clz,waw_hazard_hit {
      option.weight = 1;
   }

   //Cross CLZ instruction and RAW hazard
   cr_clz_raw_hazard: cross clz,raw_hazard_hit {
      option.weight = 1;
   }

   //CTZ instruction crosspoints
   //Cross CTZ instruction and register assignment
   cr_ctz_rs1_rd: cross ctz,rs1_addr,rd_addr {
      option.weight = 1;
   }

   //Cross CTZ instruction and RS1 toggle bits
   cr_ctz_rs1_val: cross ctz,rs1_val {
      option.weight = 1;
   }

   //Cross CTZ instruction and RS1 special values
   cr_ctz_rs1_sp_val: cross ctz,rs1_sp_val {
      option.weight = 1;
   }

   //Cross CTZ instruction and RD toggle bits
   cr_ctz_rd_val: cross ctz,rd_val {
      option.weight = 1;
   }

   //Cross CTZ instruction and RD special values
   cr_ctz_rd_sp_val: cross ctz,rd_sp_val {
      option.weight = 1;
   }

   //Cross CTZ instruction and WAR hazard
   cr_ctz_war_hazard: cross ctz,war_hazard_hit {
      option.weight = 1;
   }

   //Cross CTZ instruction and WAW hazard
   cr_ctz_waw_hazard: cross ctz,waw_hazard_hit {
      option.weight = 1;
   }

   //Cross CTZ instruction and RAW hazard
   cr_ctz_raw_hazard: cross ctz,raw_hazard_hit {
      option.weight = 1;
   }

   //CPOP instruction crosspoints
   //Cross CPOP instruction and register assignment
   cr_cpop_rs1_rd: cross cpop,rs1_addr,rd_addr {
      option.weight = 1;
   }

   //Cross CPOP instruction and RS1 toggle bits
   cr_cpop_rs1_val: cross cpop,rs1_val {
      option.weight = 1;
   }

   //Cross CPOP instruction and RS1 special values
   cr_cpop_rs1_sp_val: cross cpop,rs1_sp_val {
      option.weight = 1;
   }

   //Cross CPOP instruction and RD toggle bits
   cr_cpop_rd_val: cross cpop,rd_val {
      option.weight = 1;
   }

   //Cross CPOP instruction and RD special values
   cr_cpop_rd_sp_val: cross cpop,rd_sp_val {
      option.weight = 1;
   }

   //Cross CPOP instruction and WAR hazard
   cr_cpop_war_hazard: cross cpop,war_hazard_hit {
      option.weight = 1;
   }

   //Cross CPOP instruction and WAW hazard
   cr_cpop_waw_hazard: cross cpop,waw_hazard_hit {
      option.weight = 1;
   }

   //Cross CPOP instruction and RAW hazard
   cr_cpop_raw_hazard: cross cpop,raw_hazard_hit {
      option.weight = 1;
   }

   //MAX instruction crosspoints
   //Cross MAX instruction and register assignment
   cr_max_rs1_rs2_rd: cross max,rs1_addr,rs2_addr,rd_addr {
      option.weight = 1;
   }

   //Cross MAX instruction and RS1 toggle bits
   cr_max_rs1_val: cross max,rs1_val {
      option.weight = 1;
   }

   //Cross MAX instruction and RS1 special values
   cr_max_rs1_sp_val: cross max,rs1_sp_val {
      option.weight = 1;
   }

   //Cross MAX instruction and RS1 value sign
   cr_max_rs1_val_sign: cross max,rs1_val_sign {
      option.weight = 1;
   }

   //Cross MAX instruction and RS2 toggle bits
   cr_max_rs2_val: cross max,rs2_val {
      option.weight = 1;
   }

   //Cross MAX instruction and RS2 special values
   cr_max_rs2_sp_val: cross max,rs2_sp_val {
      option.weight = 1;
   }

   //Cross MAX instruction and RS2 value sign
   cr_max_rs2_val_sign: cross max,rs2_val_sign {
      option.weight = 1;
   }

   //Cross MAX instruction and RD toggle bits
   cr_max_rd_val: cross max,rd_val {
      option.weight = 1;
   }

   //Cross MAX instruction and RD special values
   cr_max_rd_sp_val: cross max,rd_sp_val {
      option.weight = 1;
   }

   //Cross MAX instruction and RD value sign
   cr_max_rd_val_sign: cross max,rd_val_sign {
      option.weight = 1;
   }

   //Cross MAX instruction and WAR hazard
   cr_max_war_hazard: cross max,war_hazard_hit {
      option.weight = 1;
   }

   //Cross MAX instruction and WAW hazard
   cr_max_waw_hazard: cross max,waw_hazard_hit {
      option.weight = 1;
   }

   //Cross MAX instruction and RAW hazard
   cr_max_raw_hazard: cross max,raw_hazard_hit {
      option.weight = 1;
   }

   //MAXU instruction crosspoints
   //Cross MAXU instruction and register assignment
   cr_maxu_rs1_rs2_rd: cross maxu,rs1_addr,rs2_addr,rd_addr {
      option.weight = 1;
   }

   //Cross MAXU instruction and RS1 toggle bits
   cr_maxu_rs1_val: cross maxu,rs1_val {
      option.weight = 1;
   }

   //Cross MAXU instruction and RS1 special values
   cr_maxu_rs1_sp_val: cross maxu,rs1_sp_val {
      option.weight = 1;
   }

   //Cross MAXU instruction and RS2 toggle bits
   cr_maxu_rs2_val: cross maxu,rs2_val {
      option.weight = 1;
   }

   //Cross MAXU instruction and RS2 special values
   cr_maxu_rs2_sp_val: cross maxu,rs2_sp_val {
      option.weight = 1;
   }

   //Cross MAXU instruction and RD toggle bits
   cr_maxu_rd_val: cross maxu,rd_val {
      option.weight = 1;
   }

   //Cross MAXU instruction and RD special values
   cr_maxu_rd_sp_val: cross maxu,rd_sp_val {
      option.weight = 1;
   }

   //Cross MAXU instruction and WAR hazard
   cr_maxu_war_hazard: cross maxu,war_hazard_hit {
      option.weight = 1;
   }

   //Cross MAXU instruction and WAW hazard
   cr_maxu_waw_hazard: cross maxu,waw_hazard_hit {
      option.weight = 1;
   }

   //Cross MAXU instruction and RAW hazard
   cr_maxu_raw_hazard: cross maxu,raw_hazard_hit {
      option.weight = 1;
   }

   //MIN instruction crosspoints
   //Cross MIN instruction and register assignment
   cr_min_rs1_rs2_rd: cross min,rs1_addr,rs2_addr,rd_addr {
      option.weight = 1;
   }

   //Cross MIN instruction and RS1 toggle bits
   cr_min_rs1_val: cross min,rs1_val {
      option.weight = 1;
   }

   //Cross MIN instruction and RS1 special values
   cr_min_rs1_sp_val: cross min,rs1_sp_val {
      option.weight = 1;
   }

   //Cross MIN instruction and RS1 value sign
   cr_min_rs1_val_sign: cross min,rs1_val_sign {
      option.weight = 1;
   }

   //Cross MIN instruction and RS2 toggle bits
   cr_min_rs2_val: cross min,rs2_val {
      option.weight = 1;
   }

   //Cross MIN instruction and RS2 special values
   cr_min_rs2_sp_val: cross min,rs2_sp_val {
      option.weight = 1;
   }

   //Cross MIN instruction and RS2 value sign
   cr_min_rs2_val_sign: cross min,rs2_val_sign {
      option.weight = 1;
   }

   //Cross MIN instruction and RD toggle bits
   cr_min_rd_val: cross min,rd_val {
      option.weight = 1;
   }

   //Cross MIN instruction and RD special values
   cr_min_rd_sp_val: cross min,rd_sp_val {
      option.weight = 1;
   }

   //Cross MIN instruction and RD value sign
   cr_min_rd_val_sign: cross min,rd_val_sign {
      option.weight = 1;
   }

   //Cross MIN instruction and WAR hazard
   cr_min_war_hazard: cross min,war_hazard_hit {
      option.weight = 1;
   }

   //Cross MIN instruction and WAW hazard
   cr_min_waw_hazard: cross min,waw_hazard_hit {
      option.weight = 1;
   }

   //Cross MIN instruction and RAW hazard
   cr_min_raw_hazard: cross min,raw_hazard_hit {
      option.weight = 1;
   }

   //MINU instruction crosspoints
   //Cross MINU instruction and register assignment
   cr_minu_rs1_rs2_rd: cross minu,rs1_addr,rs2_addr,rd_addr {
      option.weight = 1;
   }

   //Cross MINU instruction and RS1 toggle bits
   cr_minu_rs1_val: cross minu,rs1_val {
      option.weight = 1;
   }

   //Cross MINU instruction and RS1 special values
   cr_minu_rs1_sp_val: cross minu,rs1_sp_val {
      option.weight = 1;
   }

   //Cross MINU instruction and RS2 toggle bits
   cr_minu_rs2_val: cross minu,rs2_val {
      option.weight = 1;
   }

   //Cross MINU instruction and RS2 special values
   cr_minu_rs2_sp_val: cross minu,rs2_sp_val {
      option.weight = 1;
   }

   //Cross MINU instruction and RD toggle bits
   cr_minu_rd_val: cross minu,rd_val {
      option.weight = 1;
   }

   //Cross MINU instruction and RD special values
   cr_minu_rd_sp_val: cross minu,rd_sp_val {
      option.weight = 1;
   }

   //Cross MINU instruction and WAR hazard
   cr_minu_war_hazard: cross minu,war_hazard_hit {
      option.weight = 1;
   }

   //Cross MINU instruction and WAW hazard
   cr_minu_waw_hazard: cross minu,waw_hazard_hit {
      option.weight = 1;
   }

   //Cross MINU instruction and RAW hazard
   cr_minu_raw_hazard: cross minu,raw_hazard_hit {
      option.weight = 1;
   }

   //SEXT.B instruction crosspoints
   //Cross SEXT.B instruction and register assignment
   cr_sext_blddd_rs1__rd: cross sext_b,rs1_addr,rd_addr {
      option.weight = 1;
   }

   //Cross SEXT.B instruction and RS1 toggle bits
   cr_sext_b_rs1_val: cross sext_b,rs1_val {
      option.weight = 1;
   }

   //Cross SEXT.B instruction and RS1 special values
   cr_sext_b_rs1_sp_val: cross sext_b,rs1_sp_val {
      option.weight = 1;
   }

   //Cross SEXT.B instruction and RD toggle bits
   cr_sext_b_rd_val: cross sext_b,rd_val {
      option.weight = 1;
   }

   //Cross SEXT.B instruction and RD special values
   cr_sext_b_rd_sp_val: cross sext_b,rd_sp_val {
      option.weight = 1;
   }

   //Cross SEXT.B instruction and WAR hazard
   cr_sext_b_war_hazard: cross sext_b,war_hazard_hit {
      option.weight = 1;
   }

   //Cross SEXT.B instruction and WAW hazard
   cr_sext_b_waw_hazard: cross sext_b,waw_hazard_hit {
      option.weight = 1;
   }

   //Cross SEXT.B instruction and RAW hazard
   cr_sext_b_raw_hazard: cross sext_b,raw_hazard_hit {
      option.weight = 1;
   }

   //SEXT.H instruction crosspoints
   //Cross SEXT.H instruction and register assignment
   cr_sext_h_rs1_rd: cross sext_h,rs1_addr,rd_addr {
      option.weight = 1;
   }

   //Cross SEXT.H instruction and RS1 toggle bits
   cr_sext_h_rs1_val: cross sext_h,rs1_val {
      option.weight = 1;
   }

   //Cross SEXT.H instruction and RS1 special values
   cr_sext_h_rs1_sp_val: cross sext_h,rs1_sp_val {
      option.weight = 1;
   }

   //Cross SEXT.H instruction and RD toggle bits
   cr_sext_h_rd_val: cross sext_h,rd_val {
      option.weight = 1;
   }

   //Cross SEXT.H instruction and RD special values
   cr_sext_h_rd_sp_val: cross sext_h,rd_sp_val {
      option.weight = 1;
   }

   //Cross SEXT.H instruction and WAR hazard
   cr_sext_h_war_hazard: cross sext_h,war_hazard_hit {
      option.weight = 1;
   }

   //Cross SEXT.H instruction and WAW hazard
   cr_sext_h_waw_hazard: cross sext_h,waw_hazard_hit {
      option.weight = 1;
   }

   //Cross SEXT.H instruction and RAW hazard
   cr_sext_h_raw_hazard: cross sext_h,raw_hazard_hit {
      option.weight = 1;
   }

   //ZEXT.H instruction crosspoints
   //Cross ZEXT.H instruction and register assignment
   cr_zext_h_rs1_rd: cross zext_h,rs1_addr,rd_addr {
      option.weight = 1;
   }

   //Cross ZEXT.H instruction and RS1 toggle bits
   cr_zext_h_rs1_val: cross zext_h,rs1_val {
      option.weight = 1;
   }

   //Cross ZEXT.H instruction and RS1 special values
   cr_zext_h_rs1_sp_val: cross zext_h,rs1_sp_val {
      option.weight = 1;
   }

   //Cross ZEXT.H instruction and RD toggle bits
   cr_zext_h_rd_val: cross zext_h,rd_val {
      option.weight = 1;
   }

   //Cross ZEXT.H instruction and RD special values
   cr_zext_h_rd_sp_val: cross zext_h,rd_sp_val {
      option.weight = 1;
   }

   //Cross ZEXT.H instruction and WAR hazard
   cr_zext_h_war_hazard: cross zext_h,war_hazard_hit {
      option.weight = 1;
   }

   //Cross ZEXT.H instruction and WAW hazard
   cr_zext_h_waw_hazard: cross zext_h,waw_hazard_hit {
      option.weight = 1;
   }

   //Cross ZEXT.H instruction and RAW hazard
   cr_zext_h_raw_hazard: cross zext_h,raw_hazard_hit {
      option.weight = 1;
   }

   //ROL instruction crosspoints
   //Cross ROL instruction and register assignment
   cr_rol_rs1_rs2_rd: cross rol,rs1_addr,rs2_addr,rd_addr {
      option.weight = 1;
   }

   //Cross ROL instruction and RS1 toggle bits
   cr_rol_rs1_val: cross rol,rs1_val {
      option.weight = 1;
   }

   //Cross ROL instruction and RS1 special values
   cr_rol_rs1_sp_val: cross rol,rs1_sp_val {
      option.weight = 1;
   }

   //Cross ROL instruction and RS2 toggle bits
   cr_rol_rs2_val: cross rol,rs2_val {
      option.weight = 1;
   }

   //Cross ROL instruction and RS2 special values
   cr_rol_rs2_sp_val: cross rol,rs2_sp_val {
      option.weight = 1;
   }

   //Cross ROL instruction and RD toggle bits
   cr_rol_rd_val: cross rol,rd_val {
      option.weight = 1;
   }

   //Cross ROL instruction and RD special values
   cr_rol_rd_sp_val: cross rol,rd_sp_val {
      option.weight = 1;
   }

   //Cross ROL instruction and WAR hazard
   cr_rol_war_hazard: cross rol,war_hazard_hit {
      option.weight = 1;
   }

   //Cross ROL instruction and WAW hazard
   cr_rol_waw_hazard: cross rol,waw_hazard_hit {
      option.weight = 1;
   }

   //Cross ROL instruction and RAW hazard
   cr_rol_raw_hazard: cross rol,raw_hazard_hit {
      option.weight = 1;
   }

   //ROR instruction crosspoints
   //Cross ROR instruction and register assignment
   cr_ror_rs1_rs2_rd: cross ror,rs1_addr,rs2_addr,rd_addr {
      option.weight = 1;
   }

   //Cross ROR instruction and RS1 toggle bits
   cr_ror_rs1_val: cross ror,rs1_val {
      option.weight = 1;
   }

   //Cross ROR instruction and RS1 special values
   cr_ror_rs1_sp_val: cross ror,rs1_sp_val {
      option.weight = 1;
   }

   //Cross ROR instruction and RS2 toggle bits
   cr_ror_rs2_val: cross ror,rs2_val {
      option.weight = 1;
   }

   //Cross ROR instruction and RS2 special values
   cr_ror_rs2_sp_val: cross ror,rs2_sp_val {
      option.weight = 1;
   }

   //Cross ROR instruction and RD toggle bits
   cr_ror_rd_val: cross ror,rd_val {
      option.weight = 1;
   }

   //Cross ROR instruction and RD special values
   cr_ror_rd_sp_val: cross ror,rd_sp_val {
      option.weight = 1;
   }

   //Cross ROR instruction and WAR hazard
   cr_ror_war_hazard: cross ror,war_hazard_hit {
      option.weight = 1;
   }

   //Cross ROR instruction and WAW hazard
   cr_ror_waw_hazard: cross ror,waw_hazard_hit {
      option.weight = 1;
   }

   //Cross ROR instruction and RAW hazard
   cr_ror_raw_hazard: cross ror,raw_hazard_hit {
      option.weight = 1;
   }

   //RORI instruction crosspoints
   //Cross RORI instruction and register assignment
   cr_rori_rs1_rd: cross rori,rs1_addr,rd_addr {
      option.weight = 1;
   }

   //Cross RORI instruction and shamt toggle bits
   cr_rori_shamt_val: cross ror,shamt_val {
      option.weight = 1;
   }

   //Cross RORI instruction and shamt special values
   cr_rori_shamt_sp_val: cross rori,shamt_sp_val {
      option.weight = 1;
   }

   //Cross RORI instruction and RS1 toggle bits
   cr_rori_rs2_val: cross rori,rs1_val {
      option.weight = 1;
   }

   //Cross RORI instruction and RS1 special values
   cr_rori_rs2_sp_val: cross rori,rs1_sp_val {
      option.weight = 1;
   }

   //Cross RORI instruction and RD toggle bits
   cr_rori_rd_val: cross rori,rd_val {
      option.weight = 1;
   }

   //Cross RORI instruction and RD special values
   cr_rori_rd_sp_val: cross rori,rd_sp_val {
      option.weight = 1;
   }

   //Cross RORI instruction and WAR hazard
   cr_rori_war_hazard: cross rori,war_hazard_hit {
      option.weight = 1;
   }

   //Cross RORI instruction and WAW hazard
   cr_rori_waw_hazard: cross rori,waw_hazard_hit {
      option.weight = 1;
   }

   //Cross RORI instruction and RAW hazard
   cr_rori_raw_hazard: cross rori,raw_hazard_hit {
      option.weight = 1;
   }

   //ORC.B instruction crosspoints
   //Cross ORC.B instruction and register assignment
   cr_orc_b_rs1_rd: cross orc_b,rs1_addr,rd_addr {
      option.weight = 1;
   }

   //Cross ORC.B instruction and RS1 toggle bits
   cr_orc_b_rs1_val: cross orc_b,rs1_val {
      option.weight = 1;
   }

   //Cross ORC.B instruction and RS1 special values
   cr_orc_b_rs1_sp_val: cross orc_b,rs1_sp_val {
      option.weight = 1;
   }

   //Cross ORC.B instruction and RD toggle bits
   cr_orc_b_rd_val: cross orc_b,rd_val {
      option.weight = 1;
   }

   //Cross ORC.B instruction and RD special values
   cr_orc_b_rd_sp_val: cross orc_b,rd_sp_val {
      option.weight = 1;
   }

   //Cross ORC.B instruction and WAR hazard
   cr_orc_b_war_hazard: cross orc_b,war_hazard_hit {
      option.weight = 1;
   }

   //Cross ORC.B instruction and WAW hazard
   cr_orc_b_waw_hazard: cross orc_b,waw_hazard_hit {
      option.weight = 1;
   }

   //Cross ORC.B instruction and RAW hazard
   cr_orc_b_raw_hazard: cross orc_b,raw_hazard_hit {
      option.weight = 1;
   }

   //REV8 instruction crosspoints
   //Cross REV8 instruction and register assignment
   cr_rev8_rs1_rd: cross rev8,rs1_addr,rd_addr {
      option.weight = 1;
   }

   //Cross REV8 instruction and RS1 toggle bits
   cr_rev8_rs1_val: cross rev8,rs1_val {
      option.weight = 1;
   }

   //Cross REV8 instruction and RS1 special values
   cr_rev8_rs1_sp_val: cross rev8,rs1_sp_val {
      option.weight = 1;
   }

   //Cross REV8 instruction and RD toggle bits
   cr_rev8_rd_val: cross rev8,rd_val {
      option.weight = 1;
   }

   //Cross REV8 instruction and RD special values
   cr_rev8_rd_sp_val: cross rev8,rd_sp_val {
      option.weight = 1;
   }

   //Cross REV8 instruction and WAR hazard
   cr_rev8_war_hazard: cross rev8,war_hazard_hit {
      option.weight = 1;
   }

   //Cross REV8 instruction and WAW hazard
   cr_rev8_waw_hazard: cross rev8,waw_hazard_hit {
      option.weight = 1;
   }

   //Cross REV8 instruction and RAW hazard
   cr_rev8_raw_hazard: cross rev8,raw_hazard_hit {
      option.weight = 1;
   }

endgroup
